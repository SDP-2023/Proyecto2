module LCD_SYNC(
    input CLK, RST_n,
    output reg NCLK, GREST, HD, DEN, VD,
    output reg [11:0] Columna,
    output reg [9:0] Fila
);
    
endmodule
